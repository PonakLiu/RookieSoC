`include "include/stddef.h"
`include "chip/cpu/cpu.h"
`include "chip/cpu/isa.h"

module spm (
    
);
    
endmodule