`include "include/stddef.h"
`include "bus/bus.h"

module bus_slave_mux (
    input wire cs_0_,
    input wire cs_1_,
    input wire cs_2_,
    input wire cs_3_,
    input wire cs_4_,
    input wire cs_5_,
    input wire cs_6_,
    input wire cs_7_
);

endmodule //bus_slave_mux